// Q2: Exercise question 2.10. Provide an RTL diagram and its relevant code; also test your code using a stimulus. Keep the input and output bit size equal to 4 bits.
// y[n] = x[n] - x[n-1] + x[n-2] + x[n-3] + 0.5y[n-1] + 0.25y[n-2]

module (x,
        y);
    input x,
    output y;
    
    
endmodule

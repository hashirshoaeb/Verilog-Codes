module get_Index();
    input i, j;
    output l0,l1,l2,l3,l4,l5,l6;

    always@()
    begin
        
    end
endmodule